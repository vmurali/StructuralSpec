PrimitiveNormal.bsv