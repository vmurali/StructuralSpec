../Primitive.bsv