PrimitiveElastic.bsv