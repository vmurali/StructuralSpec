../../../lib/PrimitiveElastic.bsv