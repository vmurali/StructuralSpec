importBsv Primitive;

interface Action#(type t);
  Output#(t)
endinterface
