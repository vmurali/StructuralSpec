../../../lib/PrimitiveNormal.bsv